module graph_mem
(   
    input en,
	input clk,
	input RW,
	input data_in,
	input [4:0] coladdr,
	input [4:0] rowaddr,
	output [4:0] data_out 
);
reg [31:0] mem [31:0];
initial begin
    mem [0] = 32'b00100110001001100001011101001101;
    mem [1] = 32'b00101001010101001000100110101110;
    mem [2] = 32'b00010010100001001100101101010000;
    mem [3] = 32'b10000001110010001001100000000000;
    mem [4] = 32'b10010100010100011010100000110010;
    mem [5] = 32'b01010000010000010010010100000001;
    mem [6] = 32'b10011000000100100000000001100010;
    mem [7] = 32'b00000001000100011100001110000000;
    mem [8] = 32'b00010000100000000110000100111100;
    mem [9] = 32'b00000000000000100000010011000010;
    mem [10] = 32'b11101000001000001000000000001110;
    mem [11] = 32'b01100000110000101110101011000000;
    mem [12] = 32'b00000110010011010110000100100000;
    mem [13] = 32'b00001100000111010010001000111101;
    mem [14] = 32'b01110000000100000011010011010010;
    mem [15] = 32'b10001010010000111100010010001110;
    mem [16] = 32'b10001001010010111001100001001110;
    mem [17] = 32'b00010011101010010100100010101001;
    mem [18] = 32'b00000110000100100100100101101001;
    mem [19] = 32'b00100011010100100101010101110101;
    mem [20] = 32'b11000001001010001110100100000000;
    mem [21] = 32'b10000000000100010010000010100010;
    mem [22] = 32'b00100011001000000100100100010001;
    mem [23] = 32'b10000100000100001100010001110000;
    mem [24] = 32'b00101000000110000010000111000000;
    mem [25] = 32'b00000000101000001110100010011000;
    mem [26] = 32'b00111011100100001000000001001010;
    mem [27] = 32'b01010000010000101001101000100000;
    mem [28] = 32'b01001011111001000001111000100001;
    mem [29] = 32'b00000110001000000111100010001000;
    mem [30] = 32'b00010010100100100001000001010001;
    mem [31] = 32'b00110000010110001110000000111110;
end
reg [31:0] out_temp ;
always @ (posedge clk)begin
    if(en) begin
        if(RW) begin
        out_temp <= mem[coladdr];
        end
        else begin
           mem[coladdr][rowaddr] <= data_in;
        end
    end
    
	//data_out <= {out_temp[rowaddr+4],out_temp[rowaddr+3],out_temp[rowaddr+2],out_temp[rowaddr+1],out_temp[rowaddr]};
end
assign data_out = {out_temp[rowaddr+4],out_temp[rowaddr+3],out_temp[rowaddr+2],out_temp[rowaddr+1],out_temp[rowaddr]};
endmodule